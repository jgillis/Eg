EEN GYRATOR

Vin 1 0 5
R1 1 2 10
RC 1 3 complex(0,10)
